scan.wallpaper.walloff
scan.installs.installson
scan.startup.startoff
scan.runtime.runtimeon