scan.wallpaper.walloff
scan.installs.installsoff
scan.startup.startoff
scan.runtime.runtimeoff