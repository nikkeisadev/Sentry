127.0.0.1 cornhub.website
127.0.0.1 www.cornhub.website
