scan.wallpaper.wallon
scan.installs.installson
scan.startup.starton
scan.runtime.runtimeoff