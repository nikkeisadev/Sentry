auto_scan_mode$on
wallpaper_protection$on
runtime_check$on
directory_scan$on
installations$on
webblock$on