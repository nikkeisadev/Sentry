scan.wallpaper.wallon
scan.installs.installson
scan.startup.startoff
scan.runtime.runtimeoff